//alu.svh header file
`include "1.alu_if.sv"
`include "2.alu.sv"
`include "3.alu_tx.sv"
`include "4.alu_gen.sv"
`include "5.alu_drv.sv"
`include "6.alu_mon.sv"
`include "7.alu_scb.sv"
`include "8.alu_cov.sv"
`include "9.alu_env.sv"
`include "10.alu_tb.sv"
`include "11.alu_cfg.sv"
`include "12.alu_top.sv"
