//fifo.svh header file
`include "1.fifo_if.sv"
`include "2.fifo.sv"
`include "3.fifo_tx.sv"
`include "4.fifo_gen.sv"
`include "5.fifo_drv.sv"
`include "6.fifo_mon.sv"
`include "7.fifo_scb.sv"
`include "8.fifo_env.sv"
`include "9.fifo_tb.sv"
`include "10.fifo_cfg.sv"
`include "11.fifo_top.sv"
