`include "1.spi_if.sv"
`include "2.spi.sv"
`include "3.spi_transaction.sv"
`include "4.spi_generator.sv"
`include "5.spi_driver.sv"
`include "6.spi_monitor.sv"
`include "7.spi_scoreboard.sv"
`include "8.spi_environment.sv"
`include "9.spi_tb.sv"
`include "10.spi_cfg.sv"
