class transaction;
  
 rand bit newd;
 rand bit [11:0] din;
 bit cs;
 bit mosi;
  
  
 function void display (input string tag);
  $display("[%0s] : DATA_NEW : %0b DIN : %0d CS : %b MOSI : %0b ", tag, newd, din, cs, mosi);    
 endfunction
  
 function transaction copy();
  copy = new();
  copy.newd = this.newd;
  copy.din = this.din;
  copy.cs = this.cs;
  copy.mosi = this.mosi;
 endfunction
  
endclass
